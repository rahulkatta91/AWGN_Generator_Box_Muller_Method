
//Table with Sin/Cos Coefficient values

module Sin_Cos_Coeffs (
clk,     // Clock
address, // Address input
data    // Data output
);
input clk;
input [6:0] address;
output [30:0] data;
reg [30:0] data ;
       
always@(clk)
begin
case(address)
0 : data = 31'b 0000000011001001000_011001001000;		//Coefficient values
1 : data = 31'b 0000000011001001000_010010010000;
2 : data = 31'b 0000000011001000111_001011010111;
3 : data = 31'b 0000000011001000111_000100011100;
4 : data = 31'b 0000000011001000110_011101011110;
5 : data = 31'b 0000000011001000100_010110011101;
6 : data = 31'b 0000000011001000011_001111010111;
7 : data = 31'b 0000000011001000001_001000001101;
8 : data = 31'b 0000000011000111111_000000111110;
9 : data = 31'b 0000000011000111101_011001101000;
10 : data = 31'b 0000000011000111011_010010001011;
11 : data = 31'b 0000000011000111000_001010100110;
12 : data = 31'b 0000000011000110101_000010111001;
13 : data = 31'b 0000000011000110010_011011000100;
14 : data = 31'b 0000000011000101111_010011000100;
15 : data = 31'b 0000000011000101011_001010111001;
16 : data = 31'b 0000000011000100111_000010100100;
17 : data = 31'b 0000000011000100011_011010000011;
18 : data = 31'b 0000000011000011111_010001010100;
19 : data = 31'b 0000000011000011010_001000011001;
20 : data = 31'b 0000000011000010101_011111010000;
21 : data = 31'b 0000000011000010000_010101111000;
22 : data = 31'b 0000000011000001011_001100010000;
23 : data = 31'b 0000000011000000110_000010011001;
24 : data = 31'b 0000000011000000000_011000010001;
25 : data = 31'b 0000000010111111010_001101110111;
26 : data = 31'b 0000000010111110100_000011001100;
27 : data = 31'b 0000000010111101101_011000001110;
28 : data = 31'b 0000000010111100111_001100111100;
29 : data = 31'b 0000000010111100000_000001010110;
30 : data = 31'b 0000000010111011001_010101011100;
31 : data = 31'b 0000000010111010001_001001001100;
32 : data = 31'b 0000000010111001010_011100100111;
33 : data = 31'b 0000000010111000010_001111101011;
34 : data = 31'b 0000000010110111010_000010010111;
35 : data = 31'b 0000000010110110010_010100101100;
36 : data = 31'b 0000000010110101001_000110101000;
37 : data = 31'b 0000000010110100001_011000001100;
38 : data = 31'b 0000000010110011000_001001010101;
39 : data = 31'b 0000000010110001111_011010000101;
40 : data = 31'b 0000000010110000101_001010011001;
41 : data = 31'b 0000000010101111100_011010010011;
42 : data = 31'b 0000000010101110010_001001110000;
43 : data = 31'b 0000000010101101000_011000110000;
44 : data = 31'b 0000000010101011110_000111010100;
45 : data = 31'b 0000000010101010100_010101011010;
46 : data = 31'b 0000000010101001001_000011000001;
47 : data = 31'b 0000000010100111110_010000001010;
48 : data = 31'b 0000000010100110011_011100110100;
49 : data = 31'b 0000000010100101000_001000111110;
50 : data = 31'b 0000000010100011101_010100100111;
51 : data = 31'b 0000000010100010001_011111110000;
52 : data = 31'b 0000000010100000110_001010010111;
53 : data = 31'b 0000000010011111010_010100011101;
54 : data = 31'b 0000000010011101101_011110000000;
55 : data = 31'b 0000000010011100001_000111000001;
56 : data = 31'b 0000000010011010101_001111011110;
57 : data = 31'b 0000000010011001000_010111011000;
58 : data = 31'b 0000000010010111011_011110101101;
59 : data = 31'b 0000000010010101110_000101011110;
60 : data = 31'b 0000000010010100001_001011101010;
61 : data = 31'b 0000000010010010011_010001010001;
62 : data = 31'b 0000000010010000110_010110010010;
63 : data = 31'b 0000000010001111000_011010101100;
64 : data = 31'b 0000000010001101010_011110100000;
65 : data = 31'b 0000000010001011100_000001101110;
66 : data = 31'b 0000000010001001101_000100010011;
67 : data = 31'b 0000000010000111111_000110010010;
68 : data = 31'b 0000000010000110000_000111101000;
69 : data = 31'b 0000000010000100010_001000010101;
70 : data = 31'b 0000000010000010011_001000011010;
71 : data = 31'b 0000000010000000100_000111110110;
72 : data = 31'b 0000000001111110100_000110101001;
73 : data = 31'b 0000000001111100101_000100110010;
74 : data = 31'b 0000000001111010101_000010010010;
75 : data = 31'b 0000000001111000110_011111000111;
76 : data = 31'b 0000000001110110110_011011010001;
77 : data = 31'b 0000000001110100110_010110110001;
78 : data = 31'b 0000000001110010110_010001100111;
79 : data = 31'b 0000000001110000101_001011110001;
80 : data = 31'b 0000000001101110101_000101001111;
81 : data = 31'b 0000000001101100100_011110000010;
82 : data = 31'b 0000000001101010100_010110001010;
83 : data = 31'b 0000000001101000011_001101100101;
84 : data = 31'b 0000000001100110010_000100010101;
85 : data = 31'b 0000000001100100001_011010011000;
86 : data = 31'b 0000000001100010000_001111101110;
87 : data = 31'b 0000000001011111110_000100011001;
88 : data = 31'b 0000000001011101101_011000010110;
89 : data = 31'b 0000000001011011011_001011100111;
90 : data = 31'b 0000000001011001010_011110001011;
91 : data = 31'b 0000000001010111000_010000000010;
92 : data = 31'b 0000000001010100110_000001001100;
93 : data = 31'b 0000000001010010100_010001101001;
94 : data = 31'b 0000000001010000010_000001011001;
95 : data = 31'b 0000000001001110000_010000011011;
96 : data = 31'b 0000000001001011110_011110110001;
97 : data = 31'b 0000000001001001100_001100011001;
98 : data = 31'b 0000000001000111001_011001010100;
99 : data = 31'b 0000000001000100111_000101100010;
100 : data = 31'b 0000000001000010100_010001000010;
101 : data = 31'b 0000000001000000001_011011110110;
102 : data = 31'b 0000000000111101111_000101111100;
103 : data = 31'b 0000000000111011100_001111010101;
104 : data = 31'b 0000000000111001001_011000000010;
105 : data = 31'b 0000000000110110110_000000000001;
106 : data = 31'b 0000000000110100011_000111010100;
107 : data = 31'b 0000000000110010000_001101111010;
108 : data = 31'b 0000000000101111101_010011110011;
109 : data = 31'b 0000000000101101010_011001000000;
110 : data = 31'b 0000000000101010110_011101100001;
111 : data = 31'b 0000000000101000011_000001010110;
112 : data = 31'b 0000000000100110000_000100011111;
113 : data = 31'b 0000000000100011100_000110111100;
114 : data = 31'b 0000000000100001001_001000101101;
115 : data = 31'b 0000000000011110101_001001110011;
116 : data = 31'b 0000000000011100010_001010001110;
117 : data = 31'b 0000000000011001110_001001111110;
118 : data = 31'b 0000000000010111011_001001000100;
119 : data = 31'b 0000000000010100111_000111011111;
120 : data = 31'b 0000000000010010011_000101010000;
121 : data = 31'b 0000000000010000000_000010010111;
122 : data = 31'b 0000000000001101100_011110110101;
123 : data = 31'b 0000000000001011000_011010101001;
124 : data = 31'b 0000000000001000101_010101110101;
125 : data = 31'b 0000000000000110001_010000010111;
126 : data = 31'b 0000000000000011101_001010010010;
127 : data = 31'b 0000000000000001001_000011100101;
endcase
end

endmodule