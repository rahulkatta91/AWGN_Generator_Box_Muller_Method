
//Table with Sqrt1 Coefficient values
module Sqrt1_Coeffs (
clk,     // Clock
address, // Address input
data    // Data output
);
input clk;
input [5:0] address;
output [31:0] data;
reg [31:0] data ;
       
always@(clk)
begin
case(address)
0 : data = 32'b00000000001011010001_010000111111;
1 : data = 32'b00000000001011001011_010110101000;
2 : data = 32'b00000000001011000110_011100001011;		//Coefficient values
3 : data = 32'b00000000001011000001_000001101001;
4 : data = 32'b00000000001010111011_000111000010;
5 : data = 32'b00000000001010110110_001100010111;
6 : data = 32'b00000000001010110001_010001100110;
7 : data = 32'b00000000001010101101_010110110001;
8 : data = 32'b00000000001010101000_011011111000;
9 : data = 32'b00000000001010100011_000000111010;
10 : data = 32'b00000000001010011111_000101111000;
11 : data = 32'b00000000001010011010_001010110010;
12 : data = 32'b00000000001010010110_001111101000;
13 : data = 32'b00000000001010010010_010100011010;
14 : data = 32'b00000000001010001101_011001001001;
15 : data = 32'b00000000001010001001_011101110100;
16 : data = 32'b00000000001010000101_000010011011;
17 : data = 32'b00000000001010000001_000110111111;
18 : data = 32'b00000000001001111101_001011100000;
19 : data = 32'b00000000001001111001_001111111110;
20 : data = 32'b00000000001001110110_010100011000;
21 : data = 32'b00000000001001110010_011000101111;
22 : data = 32'b00000000001001101110_011101000100;
23 : data = 32'b00000000001001101011_000001010101;
24 : data = 32'b00000000001001100111_000101100100;
25 : data = 32'b00000000001001100100_001001110000;
26 : data = 32'b00000000001001100000_001101111001;
27 : data = 32'b00000000001001011101_010001111111;
28 : data = 32'b00000000001001011010_010110000011;
29 : data = 32'b00000000001001010111_011010000101;
30 : data = 32'b00000000001001010011_011110000100;
31 : data = 32'b00000000001001010000_000010000000;
32 : data = 32'b00000000001001001101_000101111010;
33 : data = 32'b00000000001001001010_001001110010;
34 : data = 32'b00000000001001000111_001101101000;
35 : data = 32'b00000000001001000100_010001011011;
36 : data = 32'b00000000001001000001_010101001101;
37 : data = 32'b00000000001000111110_011000111100;
38 : data = 32'b00000000001000111100_011100101001;
39 : data = 32'b00000000001000111001_000000010100;
40 : data = 32'b00000000001000110110_000011111101;
41 : data = 32'b00000000001000110011_000111100100;
42 : data = 32'b00000000001000110001_001011001010;
43 : data = 32'b00000000001000101110_001110101101;
44 : data = 32'b00000000001000101100_010010001111;
45 : data = 32'b00000000001000101001_010101101111;
46 : data = 32'b00000000001000100111_011001001101;
47 : data = 32'b00000000001000100100_011100101001;
48 : data = 32'b00000000001000100010_000000000100;
49 : data = 32'b00000000001000011111_000011011101;
50 : data = 32'b00000000001000011101_000110110100;
51 : data = 32'b00000000001000011010_001010001010;
52 : data = 32'b00000000001000011000_001101011110;
53 : data = 32'b00000000001000010110_010000110001;
54 : data = 32'b00000000001000010100_010100000010;
55 : data = 32'b00000000001000010001_010111010010;
56 : data = 32'b00000000001000001111_011010100000;
57 : data = 32'b00000000001000001101_011101101101;
58 : data = 32'b00000000001000001011_000000111001;
59 : data = 32'b00000000001000001001_000100000011;
60 : data = 32'b00000000001000000111_000111001011;
61 : data = 32'b00000000001000000101_001010010011;
62 : data = 32'b00000000001000000011_001101011001;
63 : data = 32'b00000000001000000001_010000011110;
endcase
end

endmodule
