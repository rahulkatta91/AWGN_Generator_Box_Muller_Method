
//Table with Sin/Cos Coefficient values
`timescale 1ns/1ps
module Sin_Cos_Coeffs (
address, // Address input
data    // Data output
);
input [6:0] address;
output [30:0] data;
reg [30:0] data ;
       
always@(address)
begin
case(address)
0 : data <= 31'b011001001000_0000000000000000000;
1 : data <= 31'b011001001000_0000000000000000000;
2 : data <= 31'b011001000111_0000000000000000001;	//c1,c0
3 : data <= 31'b011001000111_0000000000000000011;
4 : data <= 31'b011001000110_0000000000000000111;
5 : data <= 31'b011001000100_0000000000000001101;
6 : data <= 31'b011001000011_0000000000000010110;
7 : data <= 31'b011001000001_0000000000000100001;
8 : data <= 31'b011000111111_0000000000000110001;
9 : data <= 31'b011000111101_0000000000001000100;
10 : data <= 31'b011000111011_0000000000001011101;
11 : data <= 31'b011000111000_0000000000001111010;
12 : data <= 31'b011000110101_0000000000010011101;
13 : data <= 31'b011000110010_0000000000011000101;
14 : data <= 31'b011000101111_0000000000011110101;
15 : data <= 31'b011000101011_0000000000100101011;
16 : data <= 31'b011000100111_0000000000101101000;
17 : data <= 31'b011000100011_0000000000110101110;
18 : data <= 31'b011000011111_0000000000111111100;
19 : data <= 31'b011000011010_0000000001001010010;
20 : data <= 31'b011000010101_0000000001010110010;
21 : data <= 31'b011000010000_0000000001100011100;
22 : data <= 31'b011000001011_0000000001110010000;
23 : data <= 31'b011000000110_0000000010000001110;
24 : data <= 31'b011000000000_0000000010010011000;
25 : data <= 31'b010111111010_0000000010100101101;
26 : data <= 31'b010111110100_0000000010111001110;
27 : data <= 31'b010111101101_0000000011001111011;
28 : data <= 31'b010111100111_0000000011100110101;
29 : data <= 31'b010111100000_0000000011111111101;
30 : data <= 31'b010111011001_0000000100011010010;
31 : data <= 31'b010111010001_0000000100110110101;
32 : data <= 31'b010111001010_0000000101010100111;
33 : data <= 31'b010111000010_0000000101110100111;
34 : data <= 31'b010110111010_0000000110010110111;
35 : data <= 31'b010110110010_0000000110111010111;
36 : data <= 31'b010110101001_0000000111100000111;
37 : data <= 31'b010110100001_0000001000001000111;
38 : data <= 31'b010110011000_0000001000110011001;
39 : data <= 31'b010110001111_0000001001011111011;
40 : data <= 31'b010110000101_0000001010001101111;
41 : data <= 31'b010101111100_0000001010111110110;
42 : data <= 31'b010101110010_0000001011110001110;
43 : data <= 31'b010101101000_0000001100100111010;
44 : data <= 31'b010101011110_0000001101011111000;
45 : data <= 31'b010101010100_0000001110011001010;
46 : data <= 31'b010101001001_0000001111010110000;
47 : data <= 31'b010100111110_0000010000010101010;
48 : data <= 31'b010100110011_0000010001010111000;
49 : data <= 31'b010100101000_0000010010011011011;
50 : data <= 31'b010100011101_0000010011100010100;
51 : data <= 31'b010100010001_0000010100101100001;
52 : data <= 31'b010100000110_0000010101111000101;
53 : data <= 31'b010011111010_0000010111000111110;
54 : data <= 31'b010011101101_0000011000011001110;
55 : data <= 31'b010011100001_0000011001101110100;
56 : data <= 31'b010011010101_0000011011000110010;
57 : data <= 31'b010011001000_0000011100100000110;
58 : data <= 31'b010010111011_0000011101111110010;
59 : data <= 31'b010010101110_0000011111011110101;
60 : data <= 31'b010010100001_0000100001000010001;
61 : data <= 31'b010010010011_0000100010101000100;
62 : data <= 31'b010010000110_0000100100010010000;
63 : data <= 31'b010001111000_0000100101111110100;
64 : data <= 31'b010001101010_0000100111101110010;
65 : data <= 31'b010001011100_0000101001100001000;
66 : data <= 31'b010001001101_0000101011010111000;
67 : data <= 31'b010000111111_0000101101010000000;
68 : data <= 31'b010000110000_0000101111001100011;
69 : data <= 31'b010000100010_0000110001001011111;
70 : data <= 31'b010000010011_0000110011001110110;
71 : data <= 31'b010000000100_0000110101010100110;
72 : data <= 31'b001111110100_0000110111011110001;
73 : data <= 31'b001111100101_0000111001101010110;
74 : data <= 31'b001111010101_0000111011111010101;
75 : data <= 31'b001111000110_0000111110001101111;
76 : data <= 31'b001110110110_0001000000100100100;
77 : data <= 31'b001110100110_0001000010111110100;
78 : data <= 31'b001110010110_0001000101011011111;
79 : data <= 31'b001110000101_0001000111111100101;
80 : data <= 31'b001101110101_0001001010100000110;
81 : data <= 31'b001101100100_0001001101001000010;
82 : data <= 31'b001101010100_0001001111110011001;
83 : data <= 31'b001101000011_0001010010100001100;
84 : data <= 31'b001100110010_0001010101010011010;
85 : data <= 31'b001100100001_0001011000001000100;
86 : data <= 31'b001100010000_0001011011000001001;
87 : data <= 31'b001011111110_0001011101111101001;
88 : data <= 31'b001011101101_0001100000111100101;
89 : data <= 31'b001011011011_0001100011111111101;
90 : data <= 31'b001011001010_0001100111000101111;
91 : data <= 31'b001010111000_0001101010001111110;
92 : data <= 31'b001010100110_0001101101011100111;
93 : data <= 31'b001010010100_0001110000101101100;
94 : data <= 31'b001010000010_0001110100000001101;
95 : data <= 31'b001001110000_0001110111011001000;
96 : data <= 31'b001001011110_0001111010110011111;
97 : data <= 31'b001001001100_0001111110010010001;
98 : data <= 31'b001000111001_0010000001110011101;
99 : data <= 31'b001000100111_0010000101011000101;
100 : data <= 31'b001000010100_0010001001000001000;
101 : data <= 31'b001000000001_0010001100101100101;
102 : data <= 31'b000111101111_0010010000011011101;
103 : data <= 31'b000111011100_0010010100001101111;
104 : data <= 31'b000111001001_0010011000000011011;
105 : data <= 31'b000110110110_0010011011111100010;
106 : data <= 31'b000110100011_0010011111111000010;
107 : data <= 31'b000110010000_0010100011110111101;
108 : data <= 31'b000101111101_0010100111111010001;
109 : data <= 31'b000101101010_0010101011111111110;
110 : data <= 31'b000101010110_0010110000001000100;
111 : data <= 31'b000101000011_0010110100010100100;
112 : data <= 31'b000100110000_0010111000100011100;
113 : data <= 31'b000100011100_0010111100110101101;
114 : data <= 31'b000100001001_0011000001001010110;
115 : data <= 31'b000011110101_0011000101100010111;
116 : data <= 31'b000011100010_0011001001111110000;
117 : data <= 31'b000011001110_0011001110011100001;
118 : data <= 31'b000010111011_0011010010111101000;
119 : data <= 31'b000010100111_0011010111100000111;
120 : data <= 31'b000010010011_0011011100000111100;
121 : data <= 31'b000010000000_0011100000110001000;
122 : data <= 31'b000001101100_0011100101011101001;
123 : data <= 31'b000001011000_0011101010001100001;
124 : data <= 31'b000001000101_0011101110111101101;
125 : data <= 31'b000000110001_0011110011110001111;
126 : data <= 31'b000000011101_0011111000101000110;
127 : data <= 31'b000000001001_0011111101100010000;
endcase
end

endmodule