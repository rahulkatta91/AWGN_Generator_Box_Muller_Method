//Table with Log Coefficient values

module Log_Coeffs (
clk,     // Clock
address, // Address input
data    // Data output
);
input clk;
input [7:0] address;
output [64:0] data;
reg [64:0] data ;
       
always@(clk)
begin
case(address)
0 : data = 65'b0000000000000_1111111111000000000001_000000000000000000000000000000;
1 : data = 65'b0000000000000_1111111111111111000010_110111111000001011101100101101;
2 : data = 65'b0000000000000_0000000000111101000100_111111010001010010011011100000;
3 : data = 65'b0000000000000_0000000001111010001011_010101110100100101000011011001;		//Coefficient values
4 : data = 65'b0000000000000_0000000010110110010110_011011001011110101101010101011;
5 : data = 65'b0000000000000_0000000011110001100110_001111000001010110110000111111;
6 : data = 65'b0000000000000_0000000100101011111101_010000111111111010011011001111;
7 : data = 65'b0000000000000_0000000101100101011010_000000110010110001100000101001;
8 : data = 65'b0000000000000_0000000110011110000001_011110000101101010111001011100;
9 : data = 65'b0000000000000_0000000111010101110000_001000100100110010101110111000;
10 : data = 65'b0000000000000_0000001000001100101001_011111111100110001101100100110;
11 : data = 65'b0000000000000_0000001001000010101110_000011111010101100010011001111;
12 : data = 65'b0000000000000_0000001001110111111110_010100001100000010001100011001;
13 : data = 65'b0000000000000_0000001010101100011011_010000011110101101011111110001;
14 : data = 65'b0000000000000_0000001011100000000110_011000100001000010001001011110;
15 : data = 65'b0000000000000_0000001100010010111111_001100000001101101010001011111;
16 : data = 65'b0000000000000_0000001101000101001000_001010101111110100100100001111;
17 : data = 65'b0000000000000_0000001101110110100000_010100011010110101101100010010;
18 : data = 65'b0000000000000_0000001110100111001010_001000110010100101101101000001;
19 : data = 65'b0000000000000_0000001111010111000101_000111100111010000011110010110;
20 : data = 65'b0000000000000_0000010000000110010010_010000101001011000001001011010;
21 : data = 65'b0000000000000_0000010000110100110011_000011101001110100100110001111;
22 : data = 65'b0000000000000_0000010001100010101000_000000011001110010111010010101;
23 : data = 65'b0000000000000_0000010010001111110001_000110101010110100111000001001;
24 : data = 65'b0000000000000_0000010010111100001111_010110001110110000011111010010;
25 : data = 65'b0000000000000_0000010011101000000011_001110110111101111011101111110;
26 : data = 65'b0000000000000_0000010100010011001110_010000011000001110110010110100;
27 : data = 65'b0000000000000_0000010100111101110001_011010100010111110001111101001;
28 : data = 65'b0000000000000_0000010101100111101011_001101001010111111111101001100;
29 : data = 65'b0000000000000_0000010110010000111110_001000000011100111111111010010;
30 : data = 65'b0000000000000_0000010110111001101010_001011000000011011111001111100;
31 : data = 65'b0000000000000_0000010111100001110000_010101110101010010010111001010;
32 : data = 65'b0000000000000_0000011000001001010000_001000010110010010101101010000;
33 : data = 65'b0000000000000_0000011000110000001100_000010010111110100100110000100;
34 : data = 65'b0000000000000_0000011001010110100011_000011101110011111100110100110;
35 : data = 65'b0000000000000_0000011001111100010110_001100001111001010110111011111;
36 : data = 65'b0000000000000_0000011010100001100110_011011101110111100101101111010;
37 : data = 65'b0000000000000_0000011011000110010011_010010000011001010010101001110;
38 : data = 65'b0000000000000_0000011011101010011110_001111000001010111011000111111;
39 : data = 65'b0000000000000_0000011100001110000111_010010011111010101101111111001;
40 : data = 65'b0000000000000_0000011100110001010000_011100010011000101000110101011;
41 : data = 65'b0000000000000_0000011101010011110111_001100010010110010101100011011;
42 : data = 65'b0000000000000_0000011101110101111111_000010010100111000111110000100;
43 : data = 65'b0000000000000_0000011110010111100111_011110001111111111010011111110;
44 : data = 65'b0000000000000_0000011110111000110000_011111111010111001101110110011;
45 : data = 65'b0000000000000_0000011111011001011010_000111001100101000100101001111;
46 : data = 65'b0000000000000_0000011111111001100110_010011111100011000010010010010;
47 : data = 65'b0000000000000_0000100000011001010100_000110000001100001000011111011;
48 : data = 65'b0000000000000_0000100000111000100101_011101010011100110101010000101;
49 : data = 65'b0000000000000_0000100001010111011001_011001101010011000000110001111;
50 : data = 65'b0000000000000_0000100001110101110000_011010111101101111011011010001;
51 : data = 65'b0000000000000_0000100010010011101100_000001000101110001011101101100;
52 : data = 65'b0000000000000_0000100010110001001100_001011111010101101100100100001;
53 : data = 65'b0000000000000_0000100011001110010001_011011010100111101011010000111;
54 : data = 65'b0000000000000_0000100011101010111011_001111001101000100101101101111;
55 : data = 65'b0000000000000_0000100100000111001011_000111011011110001000101100110;
56 : data = 65'b0000000000000_0000100100100011000001_000011111001111001110000000001;
57 : data = 65'b0000000000000_0000100100111110011101_000100100000011111010111010010;
58 : data = 65'b0000000000000_0000100101011001100001_001001001000101011110011011010;
59 : data = 65'b0000000000000_0000100101110100001011_010001101011110001111101101000;
60 : data = 65'b0000000000000_0000100110001110011101_011110000011001101100011101110;
61 : data = 65'b0000000000000_0000100110101000010111_001110001000100010111011110111;
62 : data = 65'b0000000000000_0000100111000001111001_000001110101011110111000100000;
63 : data = 65'b0000000000000_0000100111011011000011_011001000011110110011100110111;
64 : data = 65'b0000000000000_0000100111110011110111_010011101101100110110001001110;
65 : data = 65'b0000000000000_0000101000001100010100_010001101100110100111000000011;
66 : data = 65'b0000000000000_0000101000100100011010_010010111011101101100010111110;
67 : data = 65'b0000000000000_0000101000111100001010_010111010100100101001000010110;
68 : data = 65'b0000000000000_0000101001010011100101_011110110001110111011000100011;
69 : data = 65'b0000000000000_0000101001101010101010_001001001110000111010100001100;
70 : data = 65'b0000000000000_0000101010000001011010_010110100011111111000001111011;
71 : data = 65'b0000000000000_0000101010010111110101_000110101110001111100101010100;
72 : data = 65'b0000000000000_0000101010101101111100_011001100111110000110100011010;
73 : data = 65'b0000000000000_0000101011000011101110_001111001011100001001111100110;
74 : data = 65'b0000000000000_0000101011011001001101_000111010100100101111000111111;
75 : data = 65'b0000000000000_0000101011101110011000_000001111110001010001000010111;
76 : data = 65'b0000000000000_0000101100000011001111_011111000011011111100111101100;
77 : data = 65'b0000000000000_0000101100010111110011_011110011111111110000110100101;
78 : data = 65'b0000000000000_0000101100101100000101_000000001111000011010100000110;
79 : data = 65'b0000000000000_0000101101000000000100_000100001100010010110110000100;
80 : data = 65'b0000000000000_0000101101010011110000_001010010011010110000001011000;
81 : data = 65'b0000000000000_0000101101100111001011_010010011111111011110010101100;
82 : data = 65'b0000000000000_0000101101111010010100_011100101101111000100110001011;
83 : data = 65'b0000000000000_0000101110001101001011_001000111001000110010001001101;
84 : data = 65'b0000000000000_0000101110011111110001_010110111101100011111010010010;
85 : data = 65'b0000000000000_0000101110110010000101_000110110111010101110010011011;
86 : data = 65'b0000000000000_0000101111000100001001_011000100010100101010000000000;
87 : data = 65'b0000000000000_0000101111010101111101_001011111011100000100011001010;
88 : data = 65'b0000000000000_0000101111100111100000_000000111110011010110101110000;
89 : data = 65'b0000000000000_0000101111111000110010_010111100111101100000000101011;
90 : data = 65'b0000000000000_0000110000001001110101_001111110011110000100110100110;
91 : data = 65'b0000000000000_0000110000011010101000_001001011111001001101110101011;
92 : data = 65'b0000000000000_0000110000101011001100_000100100110011100111101000011;
93 : data = 65'b0000000000000_0000110000111011100001_000001000110010100001111100110;
94 : data = 65'b0000000000000_0000110001001011100110_011110111011011101110100100111;
95 : data = 65'b0000000000000_0000110001011011011100_011110000010101100001001001010;
96 : data = 65'b0000000000000_0000110001101011000100_011110011000110101110000100000;
97 : data = 65'b0000000000000_0000110001111010011101_011111111010110101010000100101;
98 : data = 65'b0000000000000_0000110010001001101001_000010100101101001001011110100;
99 : data = 65'b0000000000000_0000110010011000100110_000110010110010011111101010001;
100 : data = 65'b0000000000000_0000110010100111010101_001011001001111011110001101011;
101 : data = 65'b0000000000000_0000110010110101110110_010000111101101010100100101001;
102 : data = 65'b0000000000000_0000110011000100001010_010111101110101101111010101101;
103 : data = 65'b0000000000000_0000110011010010010001_011111011010010110111100110100;
104 : data = 65'b0000000000000_0000110011100000001010_000111111101111010010100000000;
105 : data = 65'b0000000000000_0000110011101101110110_010001010110110000000100010001;
106 : data = 65'b0000000000000_0000110011111011010110_011011100010010011101011001110;
107 : data = 65'b0000000000000_0000110100001000101001_000110011110000011110100101000;
108 : data = 65'b0000000000000_0000110100010101110000_010010000111100010011111101101;
109 : data = 65'b0000000000000_0000110100100010101010_011110011100010100110011011111;
110 : data = 65'b0000000000000_0000110100101111011000_001011011010000010111110000100;
111 : data = 65'b0000000000000_0000110100111011111010_011000111110011000010001110111;
112 : data = 65'b0000000000000_0000110101001000010001_000111000111000010111101101011;
113 : data = 65'b0000000000000_0000110101010100011011_010101110001110100001100011110;
114 : data = 65'b0000000000000_0000110101100000011010_000100111100100000000001011000;
115 : data = 65'b0000000000000_0000110101101100001110_010100100100111101010010001011;
116 : data = 65'b0000000000000_0000110101110111110111_000100101001000101100101101001;
117 : data = 65'b0000000000000_0000110110000011010100_010101000110110101001110011101;
118 : data = 65'b0000000000000_0000110110001110100111_000101111100001011001011101111;
119 : data = 65'b0000000000000_0000110110011001101111_010111000111001000111100111001;
120 : data = 65'b0000000000000_0000110110100100101100_001000100101110010101010110011;
121 : data = 65'b0000000000000_0000110110101111011111_011010010110001110111010010111;
122 : data = 65'b0000000000000_0000110110111010000111_001100010110100110101101011000;
123 : data = 65'b0000000000000_0000110111000100100101_011110100101000101100000110110;
124 : data = 65'b0000000000000_0000110111001110111001_010000111111111001000111000011;
125 : data = 65'b0000000000000_0000110111011001000100_000011100101010001100101110010;
126 : data = 65'b0000000000000_0000110111100011000100_010110010011100001010110000000;
127 : data = 65'b0000000000000_0000110111101100111010_001001001000111100111011010110;
128 : data = 65'b0000000000000_0000110111110110100111_011100000011111011000111101000;
129 : data = 65'b0000000000000_0000111000000000001011_001111000010110100110100101000;
130 : data = 65'b0000000000000_0000111000001001100101_000010000100000101000001001101;
131 : data = 65'b0000000000000_0000111000010010110110_010101000110001000110000110100;
132 : data = 65'b0000000000000_0000111000011011111110_001000000111011111000111010001;
133 : data = 65'b0000000000000_0000111000100100111101_011011000110101001000111011000;
134 : data = 65'b0000000000000_0000111000101101110011_001110000010001001110000000101;
135 : data = 65'b0000000000000_0000111000110110100000_000000111000100101111001000101;
136 : data = 65'b0000000000000_0000111000111111000101_010011101000100100010010011111;
137 : data = 65'b0000000000000_0000111001000111100001_000110010000101101100001111000;
138 : data = 65'b0000000000000_0000111001001111110101_011000101111101011111110001100;
139 : data = 65'b0000000000000_0000111001011000000000_001011000100001011101111100011;
140 : data = 65'b0000000000000_0000111001100000000011_011101001100111010110000111000;
141 : data = 65'b0000000000000_0000111001100111111110_001111001000101000100000001100;
142 : data = 65'b0000000000000_0000111001101111110001_000000110110000110001111011001;
143 : data = 65'b0000000000000_0000111001110111011100_010010010100000110110100100001;
144 : data = 65'b0000000000000_0000111001111110111111_000011100001011110101100011101;
145 : data = 65'b0000000000000_0000111010000110011011_010100011101000011110111011011;
146 : data = 65'b0000000000000_0000111010001101101111_000101000101101101111100110100;
147 : data = 65'b0000000000000_0000111010010100111100_010101011010010101111101110100;
148 : data = 65'b0000000000000_0000111010011100000001_000101011001110110100010110010;
149 : data = 65'b0000000000000_0000111010100010111110_010101000011001011101000011100;
150 : data = 65'b0000000000000_0000111010101001110101_000100010101010010101110110010;
151 : data = 65'b0000000000000_0000111010110000100100_010011001111001010101001111100;
152 : data = 65'b0000000000000_0000111010110111001100_000001101111110011101010000001;
153 : data = 65'b0000000000000_0000111010111101101110_001111110110001111010011010111;
154 : data = 65'b0000000000000_0000111011000100001000_011101100001100000011110100101;
155 : data = 65'b0000000000000_0000111011001010011100_001010110000101011011001111010;
156 : data = 65'b0000000000000_0000111011010000101000_010111100010110101100010101011;
157 : data = 65'b0000000000000_0000111011010110101111_000011110111000101101001000010;
158 : data = 65'b0000000000000_0000111011011100101110_001111101100100011101000000111;
159 : data = 65'b0000000000000_0000111011100010101000_011011000010011000101011111000;
160 : data = 65'b0000000000000_0000111011101000011010_000101110111101111001010010111;
161 : data = 65'b0000000000000_0000111011101110000111_010000001011110010100011011100;
162 : data = 65'b0000000000000_0000111011110011101101_011001111101101111100001000111;
163 : data = 65'b0000000000000_0000111011111001001101_000011001100110011110100110010;
164 : data = 65'b0000000000000_0000111011111110100111_001011111000001110010100011110;
165 : data = 65'b0000000000000_0000111100000011111011_010011111111001110111110100001;
166 : data = 65'b0000000000000_0000111100001001001001_011011100001000110110000101110;
167 : data = 65'b0000000000000_0000111100001110010010_000010011101000111110000110111;
168 : data = 65'b0000000000000_0000111100010011010100_001000110010100100111111000111;
169 : data = 65'b0000000000000_0000111100011000010001_001110100000110010100001010011;
170 : data = 65'b0000000000000_0000111100011101001000_010011100111000101011010001000;
171 : data = 65'b0000000000000_0000111100100001111001_011000000100110011101000011010;
172 : data = 65'b0000000000000_0000111100100110100101_011011111001010100001100100101;
173 : data = 65'b0000000000000_0000111100101011001100_011111000011111110111010000010;
174 : data = 65'b0000000000000_0000111100101111101101_000001100100001100100111011100;
175 : data = 65'b0000000000000_0000111100110100001001_000011011001010110111110011100;
176 : data = 65'b0000000000000_0000111100111000011111_000100100010111000100100010010;
177 : data = 65'b0000000000000_0000111100111100110001_000101000000001100110101110110;
178 : data = 65'b0000000000000_0000111101000000111101_000100110000110000000000100100;
179 : data = 65'b0000000000000_0000111101000101000100_000011110011111111001101010111;
180 : data = 65'b0000000000000_0000111101001001000110_000010001001011000011101000111;
181 : data = 65'b0000000000000_0000111101001101000011_011111110000011010010010001111;
182 : data = 65'b0000000000000_0000111101010000111100_011100101000100100010101011001;
183 : data = 65'b0000000000000_0000111101010100101111_011000110001010110110111100110;
184 : data = 65'b0000000000000_0000111101011000011110_010100001010010010111001111100;
185 : data = 65'b0000000000000_0000111101011100001000_001110110010111010001110100101;
186 : data = 65'b0000000000000_0000111101011111101101_001000101010101111010110111111;
187 : data = 65'b0000000000000_0000111101100011001110_000001110001010101100001011111;
188 : data = 65'b0000000000000_0000111101100110101010_011010000110010000101000110110;
189 : data = 65'b0000000000000_0000111101101010000010_010001101001000101011000001111;
190 : data = 65'b0000000000000_0000111101101101010101_001000011001011000111101110010;
191 : data = 65'b0000000000000_0000111101110000100100_011110010110110001011100001001;
192 : data = 65'b0000000000000_0000111101110011101110_010011100000110101011001101111;
193 : data = 65'b0000000000000_0000111101110110110101_000111110111001100000110010100;
194 : data = 65'b0000000000000_0000111101111001110111_011011011001011101011011101101;
195 : data = 65'b0000000000000_0000111101111100110101_001110000111010001111100110110;
196 : data = 65'b0000000000000_0000111101111111101110_000000000000010010101100111110;
197 : data = 65'b0000000000000_0000111110000010100100_010001000100001001011110110101;
198 : data = 65'b0000000000000_0000111110000101010110_000001010010100000100010111010;
199 : data = 65'b0000000000000_0000111110001000000011_010000101011000010110001101001;
200 : data = 65'b0000000000000_0000111110001010101101_011111001101011011100111101101;
201 : data = 65'b0000000000000_0000111110001101010011_001100111001010111000111000001;
202 : data = 65'b0000000000000_0000111110001111110101_011001101110100001101100110101;
203 : data = 65'b0000000000000_0000111110010010010011_000101101100101000100001110111;
204 : data = 65'b0000000000000_0000111110010100101101_010000110011011001001111011011;
205 : data = 65'b0000000000000_0000111110010111000100_011011000010100001110101001100;
206 : data = 65'b0000000000000_0000111110011001010111_000100011001110000111110010111;
207 : data = 65'b0000000000000_0000111110011011100110_001100111000110101110100111101;
208 : data = 65'b0000000000000_0000111110011101110010_010100011111011111111011010101;
209 : data = 65'b0000000000000_0000111110011111111010_011011001101011111011010100011;
210 : data = 65'b0000000000000_0000111110100001111111_000001000010100100110001011110;
211 : data = 65'b0000000000000_0000111110100100000000_000101111110100001000011000010;
212 : data = 65'b0000000000000_0000111110100101111110_001010000001000101110010001010;
213 : data = 65'b0000000000000_0000111110100111111001_001101001010000100101110001111;
214 : data = 65'b0000000000000_0000111110101001110000_001111011001010000010110011000;
215 : data = 65'b0000000000000_0000111110101011100100_010000101110011011010101011001;
216 : data = 65'b0000000000000_0000111110101101010100_010001001001011001000000001000;
217 : data = 65'b0000000000000_0000111110101111000010_010000101001111100110100000000;
218 : data = 65'b0000000000000_0000111110110000101100_001111001111111010111000101001;
219 : data = 65'b0000000000000_0000111110110010010011_001100111011000111100101011111;
220 : data = 65'b0000000000000_0000111110110011110111_001001101011010111101110101111;
221 : data = 65'b0000000000000_0000111110110101011000_000101100000100000011111010111;
222 : data = 65'b0000000000000_0000111110110110110110_000000011010010111011011000001;
223 : data = 65'b0000000000000_0000111110111000010000_011010011000110010011111111001;
224 : data = 65'b0000000000000_0000111110111001101000_010011011011100111111101010010;
225 : data = 65'b0000000000000_0000111110111010111101_001011100010101110011101100101;
226 : data = 65'b0000000000000_0000111110111100001111_000010101101111101000100111010;
227 : data = 65'b0000000000000_0000111110111101011110_011000111101001011000010010101;
228 : data = 65'b0000000000000_0000111110111110101011_001110010000010000000111001010;
229 : data = 65'b0000000000000_0000111110111111110100_000010100111000100010000101010;
230 : data = 65'b0000000000000_0000111111000000111011_010110000001011111110111111100;
231 : data = 65'b0000000000000_0000111111000001111111_001000011111011011100000110110;
232 : data = 65'b0000000000000_0000111111000011000000_011010000000110000010000010100;
233 : data = 65'b0000000000000_0000111111000011111111_001010100101010111010011001001;
234 : data = 65'b0000000000000_0000111111000100111011_011010001101001010001111111110;
235 : data = 65'b0000000000000_0000111111000101110100_001000111000000010111100111011;
236 : data = 65'b0000000000000_0000111111000110101011_010110100101111011101010011100;
237 : data = 65'b0000000000000_0000111111000111011111_000011010110101110101100111001;
238 : data = 65'b0000000000000_0000111111001000010001_001111001010010110110110010110;
239 : data = 65'b0000000000000_0000111111001001000000_011010000000101111001000110000;
240 : data = 65'b0000000000000_0000111111001001101101_000011111001110010110011111001;
241 : data = 65'b0000000000000_0000111111001010010111_001100110101011101011001011110;
242 : data = 65'b0000000000000_0000111111001010111111_010100110011101010101101001011;
243 : data = 65'b0000000000000_0000111111001011100101_011011110100010110110011001001;
244 : data = 65'b0000000000000_0000111111001100001000_000001110111011110000000000000;
245 : data = 65'b0000000000000_0000111111001100101001_000110111100111100110001010100;
246 : data = 65'b0000000000000_0000111111001101000111_001011000100101111111110001000;
247 : data = 65'b0000000000000_0000111111001101100011_001110001110110100100111100110;
248 : data = 65'b0000000000000_0000111111001101111101_010000011011000111111011011101;
249 : data = 65'b0000000000000_0000111111001110010101_010001101001100111011100111010;
250 : data = 65'b0000000000000_0000111111001110101011_010001111010010000110101100001;
251 : data = 65'b0000000000000_0000111111001110111110_010001001101000010000010011100;
252 : data = 65'b0000000000000_0000111111001111010000_001111100001111001001100010100;
253 : data = 65'b0000000000000_0000111111001111011111_001100111000110100101001100110;
254 : data = 65'b0000000000000_0000111111001111101100_001001010001110010111111100101;
255 : data = 65'b0000000000000_0000111111001111110111_000100101100110010111100011000;
endcase
end

endmodule
