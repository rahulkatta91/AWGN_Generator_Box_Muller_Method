
//Table with Sqrt1 Coefficient values
`timescale 1ns/1ps
module Sqrt1_Coeffs (
address, // Address input
data    // Data output
);
input [5:0] address;
output [31:0] data;
reg [31:0] data ;
       
always@(address)
begin
case(address)
0 : data <= 32'b000101101000_00101101011011100010;
1 : data <= 32'b000101100101_00101101110001111111;	//Coefficients c1,c0
2 : data <= 32'b000101100011_00101110001000010001;
3 : data <= 32'b000101100000_00101110011110011000;
4 : data <= 32'b000101011101_00101110110100010101;
5 : data <= 32'b000101011011_00101111001010001000;
6 : data <= 32'b000101011000_00101111011111110001;
7 : data <= 32'b000101010110_00101111110101010000;
8 : data <= 32'b000101010100_00110000001010100101;
9 : data <= 32'b000101010001_00110000011111110001;
10 : data <= 32'b000101001111_00110000110100110100;
11 : data <= 32'b000101001101_00110001001001101110;
12 : data <= 32'b000101001011_00110001011110011111;
13 : data <= 32'b000101001001_00110001110011000111;
14 : data <= 32'b000101000110_00110010000111100111;
15 : data <= 32'b000101000100_00110010011011111111;
16 : data <= 32'b000101000010_00110010110000001110;
17 : data <= 32'b000101000000_00110011000100010101;
18 : data <= 32'b000100111110_00110011011000010101;
19 : data <= 32'b000100111100_00110011101100001101;
20 : data <= 32'b000100111011_00110011111111111101;
21 : data <= 32'b000100111001_00110100010011100101;
22 : data <= 32'b000100110111_00110100100111000111;
23 : data <= 32'b000100110101_00110100111010100001;
24 : data <= 32'b000100110011_00110101001101110100;
25 : data <= 32'b000100110010_00110101100001000000;
26 : data <= 32'b000100110000_00110101110100000101;
27 : data <= 32'b000100101110_00110110000111000100;
28 : data <= 32'b000100101101_00110110011001111100;
29 : data <= 32'b000100101011_00110110101100101101;
30 : data <= 32'b000100101001_00110110111111011000;
31 : data <= 32'b000100101000_00110111010001111101;
32 : data <= 32'b000100100110_00110111100100011011;
33 : data <= 32'b000100100101_00110111110110110011;
34 : data <= 32'b000100100011_00111000001001000110;
35 : data <= 32'b000100100010_00111000011011010010;
36 : data <= 32'b000100100000_00111000101101011001;
37 : data <= 32'b000100011111_00111000111111011001;
38 : data <= 32'b000100011110_00111001010001010101;
39 : data <= 32'b000100011100_00111001100011001010;
40 : data <= 32'b000100011011_00111001110100111010;
41 : data <= 32'b000100011001_00111010000110100101;
42 : data <= 32'b000100011000_00111010011000001010;
43 : data <= 32'b000100010111_00111010101001101010;
44 : data <= 32'b000100010110_00111010111011000101;
45 : data <= 32'b000100010100_00111011001100011011;
46 : data <= 32'b000100010011_00111011011101101011;
47 : data <= 32'b000100010010_00111011101110110111;
48 : data <= 32'b000100010001_00111011111111111110;
49 : data <= 32'b000100001111_00111100010001000000;
50 : data <= 32'b000100001110_00111100100001111101;
51 : data <= 32'b000100001101_00111100110010110101;
52 : data <= 32'b000100001100_00111101000011101001;
53 : data <= 32'b000100001011_00111101010100011000;
54 : data <= 32'b000100001010_00111101100101000010;
55 : data <= 32'b000100001000_00111101110101101000;
56 : data <= 32'b000100000111_00111110000110001010;
57 : data <= 32'b000100000110_00111110010110100111;
58 : data <= 32'b000100000101_00111110100111000000;
59 : data <= 32'b000100000100_00111110110111010101;
60 : data <= 32'b000100000011_00111111000111100101;
61 : data <= 32'b000100000010_00111111010111110001;
62 : data <= 32'b000100000001_00111111100111111001;
63 : data <= 32'b000100000000_00111111110111111101;
endcase
end

endmodule
