//Table with Sqrt2 Coefficient values
`timescale 1ns/1ps
module Sqrt2_Coeffs (
address, // Address input
data    // Data output
);
input [5:0] address;
output [31:0] data;
reg [31:0] data ;
       
always@(address)
begin
case(address)
0 : data <= 32'b000111111110_00100000000111111100;	//c1,c0 Coefficients
1 : data <= 32'b000111111010_00100000010111110100;
2 : data <= 32'b000111110110_00100000100111100100;
3 : data <= 32'b000111110010_00100000110111001101;
4 : data <= 32'b000111101110_00100001000110101111;
5 : data <= 32'b000111101011_00100001010110001001;
6 : data <= 32'b000111100111_00100001100101011100;
7 : data <= 32'b000111100100_00100001110100101000;
8 : data <= 32'b000111100001_00100010000011101110;
9 : data <= 32'b000111011101_00100010010010101101;
10 : data <= 32'b000111011010_00100010100001100101;
11 : data <= 32'b000111010111_00100010110000010111;
12 : data <= 32'b000111010100_00100010111111000011;
13 : data <= 32'b000111010001_00100011001101101000;
14 : data <= 32'b000111001110_00100011011100001000;
15 : data <= 32'b000111001011_00100011101010100010;
16 : data <= 32'b000111001000_00100011111000110110;
17 : data <= 32'b000111000101_00100100000111000100;
18 : data <= 32'b000111000010_00100100010101001101;
19 : data <= 32'b000111000000_00100100100011010000;
20 : data <= 32'b000110111101_00100100110001001110;
21 : data <= 32'b000110111010_00100100111111000110;
22 : data <= 32'b000110111000_00100101001100111010;
23 : data <= 32'b000110110101_00100101011010101000;
24 : data <= 32'b000110110011_00100101101000010001;
25 : data <= 32'b000110110000_00100101110101110110;
26 : data <= 32'b000110101110_00100110000011010101;
27 : data <= 32'b000110101100_00100110010000110000;
28 : data <= 32'b000110101001_00100110011110000110;
29 : data <= 32'b000110100111_00100110101011011000;
30 : data <= 32'b000110100101_00100110111000100101;
31 : data <= 32'b000110100011_00100111000101101101;
32 : data <= 32'b000110100000_00100111010010110001;
33 : data <= 32'b000110011110_00100111011111110001;
34 : data <= 32'b000110011100_00100111101100101100;
35 : data <= 32'b000110011010_00100111111001100100;
36 : data <= 32'b000110011000_00101000000110010111;
37 : data <= 32'b000110010110_00101000010011000110;
38 : data <= 32'b000110010100_00101000011111110001;
39 : data <= 32'b000110010010_00101000101100011001;
40 : data <= 32'b000110010000_00101000111000111100;
41 : data <= 32'b000110001110_00101001000101011011;
42 : data <= 32'b000110001100_00101001010001110111;
43 : data <= 32'b000110001011_00101001011110001111;
44 : data <= 32'b000110001001_00101001101010100011;
45 : data <= 32'b000110000111_00101001110110110100;
46 : data <= 32'b000110000101_00101010000011000001;
47 : data <= 32'b000110000011_00101010001111001011;
48 : data <= 32'b000110000010_00101010011011010001;
49 : data <= 32'b000110000000_00101010100111010011;
50 : data <= 32'b000101111110_00101010110011010011;
51 : data <= 32'b000101111101_00101010111111001111;
52 : data <= 32'b000101111011_00101011001011000111;
53 : data <= 32'b000101111001_00101011010110111101;
54 : data <= 32'b000101111000_00101011100010101111;
55 : data <= 32'b000101110110_00101011101110011110;
56 : data <= 32'b000101110101_00101011111010001010;
57 : data <= 32'b000101110011_00101100000101110010;
58 : data <= 32'b000101110010_00101100010001011000;
59 : data <= 32'b000101110000_00101100011100111011;
60 : data <= 32'b000101101111_00101100101000011010;
61 : data <= 32'b000101101101_00101100110011110111;
62 : data <= 32'b000101101100_00101100111111010001;
63 : data <= 32'b000101101010_00101101001010101000;
endcase
end

endmodule
