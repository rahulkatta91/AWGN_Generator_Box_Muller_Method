//Table with Log Coefficient values
`timescale 1ns/1ps
module Log_Coeffs (
address, // Address input
data    // Data output
);

input [7:0] address;
output [64:0] data;
reg [64:0] data ;
       
always@(address)
begin
case(address)
0 : data <= 65'b0001111111000_1000000001111110110100_010111111100000010000100001011;	//c2,c1,c0
1 : data <= 65'b0001111110000_1000000011111100110110_010111111000000100100010010100;
2 : data <= 65'b0001111101000_1000000101111001111010_010111110100000111111111000000;
3 : data <= 65'b0001111100000_1000000111110110000000_010111110000001100011001101110;
4 : data <= 65'b0001111011001_1000001001110001001010_010111101100010001110010000010;
5 : data <= 65'b0001111010001_1000001011101011011000_010111101000011000000111011100;
6 : data <= 65'b0001111001010_1000001101100100101011_010111100100011111011001011111;
7 : data <= 65'b0001111000011_1000001111011101000011_010111100000100111100111101110;
8 : data <= 65'b0001110111011_1000010001010100100001_010111011100110000110001101100;
9 : data <= 65'b0001110110100_1000010011001011000110_010111011000111010110110111100;
10 : data <= 65'b0001110101101_1000010101000000110010_010111010101000101110111000001;
11 : data <= 65'b0001110100110_1000010110110101100110_010111010001010001110001100000;
12 : data <= 65'b0001110011111_1000011000101001100011_010111001101011110100101111101;
13 : data <= 65'b0001110011000_1000011010011100101001_010111001001101100010011111101;
14 : data <= 65'b0001110010010_1000011100001110111001_010111000101111010111011000011;
15 : data <= 65'b0001110001011_1000011110000000010011_010111000010001010011010110111;
16 : data <= 65'b0001110000100_1000011111110000111001_010110111110011010110010111100;
17 : data <= 65'b0001101111110_1000100001100000101010_010110111010101100000010111000;
18 : data <= 65'b0001101110111_1000100011001111100111_010110110110111110001010010011;
19 : data <= 65'b0001101110001_1000100100111101110001_010110110011010001001000110010;
20 : data <= 65'b0001101101011_1000100110101011001000_010110101111100100111101111011;
21 : data <= 65'b0001101100100_1000101000010111101101_010110101011111001101001010110;
22 : data <= 65'b0001101011110_1000101010000011100000_010110101000001111001010101001;
23 : data <= 65'b0001101011000_1000101011101110100011_010110100100100101100001011101;
24 : data <= 65'b0001101010010_1000101101011000110100_010110100000111100101101011001;
25 : data <= 65'b0001101001100_1000101111000010010110_010110011101010100101110000100;
26 : data <= 65'b0001101000110_1000110000101011001000_010110011001101101100011000111;
27 : data <= 65'b0001101000000_1000110010010011001011_010110010110000111001100001010;
28 : data <= 65'b0001100111010_1000110011111010011111_010110010010100001101000110110;
29 : data <= 65'b0001100110101_1000110101100001000101_010110001110111100111000110100;
30 : data <= 65'b0001100101111_1000110111000110111110_010110001011011000111011101110;
31 : data <= 65'b0001100101001_1000111000101100001010_010110000111110101110001001100;
32 : data <= 65'b0001100100100_1000111010010000101001_010110000100010011011000111000;
33 : data <= 65'b0001100011110_1000111011110100011011_010110000000110001110010011100;
34 : data <= 65'b0001100011001_1000111101010111100010_010101111101010000111101100010;
35 : data <= 65'b0001100010011_1000111110111001111110_010101111001110000111001110100;
36 : data <= 65'b0001100001110_1001000000011011101111_010101110110010001100110111110;
37 : data <= 65'b0001100001001_1001000001111100110101_010101110010110011000100101001;
38 : data <= 65'b0001100000011_1001000011011101010010_010101101111010101010010100001;
39 : data <= 65'b0001011111110_1001000100111101000101_010101101011111000010000010001;
40 : data <= 65'b0001011111001_1001000110011100001110_010101101000011011111101100100;
41 : data <= 65'b0001011110100_1001000111111010101111_010101100101000000011010000110;
42 : data <= 65'b0001011101111_1001001001011000101000_010101100001100101100101100011;
43 : data <= 65'b0001011101010_1001001010110101111001_010101011110001011011111100111;
44 : data <= 65'b0001011100101_1001001100010010100010_010101011010110010000111111101;
45 : data <= 65'b0001011100000_1001001101101110100100_010101010111011001011110010011;
46 : data <= 65'b0001011011011_1001001111001001111111_010101010100000001100010010101;
47 : data <= 65'b0001011010111_1001010000100100110100_010101010000101010010011110000;
48 : data <= 65'b0001011010010_1001010001111111000011_010101001101010011110010010000;
49 : data <= 65'b0001011001101_1001010011011000101100_010101001001111101111101100100;
50 : data <= 65'b0001011001000_1001010100110001110001_010101000110101000110101010111;
51 : data <= 65'b0001011000100_1001010110001010010000_010101000011010100011001011001;
52 : data <= 65'b0001010111111_1001010111100010001010_010101000000000000101001010110;
53 : data <= 65'b0001010111011_1001011000111001100001_010100111100101101100100111100;
54 : data <= 65'b0001010110110_1001011010010000010011_010100111001011011001011111010;
55 : data <= 65'b0001010110010_1001011011100110100010_010100110110001001011101111101;
56 : data <= 65'b0001010101101_1001011100111100001110_010100110010111000011010110101;
57 : data <= 65'b0001010101001_1001011110010001011000_010100101111101000000010001111;
58 : data <= 65'b0001010100101_1001011111100101111110_010100101100011000010011111011;
59 : data <= 65'b0001010100001_1001100000111010000011_010100101001001001001111100111;
60 : data <= 65'b0001010011100_1001100010001101100101_010100100101111010110101000011;
61 : data <= 65'b0001010011000_1001100011100000100111_010100100010101101000011111101;
62 : data <= 65'b0001010010100_1001100100110011000110_010100011111011111111100000101;
63 : data <= 65'b0001010010000_1001100110000101000101_010100011100010011011101001011;
64 : data <= 65'b0001010001100_1001100111010110100100_010100011001000111100110111110;
65 : data <= 65'b0001010001000_1001101000100111100010_010100010101111100011001001110;
66 : data <= 65'b0001010000100_1001101001111000000000_010100010010110001110011101011;
67 : data <= 65'b0001010000000_1001101011000111111111_010100001111100111110110000101;
68 : data <= 65'b0001001111100_1001101100010111011110_010100001100011110100000001101;
69 : data <= 65'b0001001111000_1001101101100110011110_010100001001010101110001110010;
70 : data <= 65'b0001001110100_1001101110110100111111_010100000110001101101010100111;
71 : data <= 65'b0001001110000_1001110000000011000001_010100000011000110001010011010;
72 : data <= 65'b0001001101101_1001110001010000100110_010011111111111111010000111110;
73 : data <= 65'b0001001101001_1001110010011101101100_010011111100111000111110000010;
74 : data <= 65'b0001001100101_1001110011101010010101_010011111001110011010001011001;
75 : data <= 65'b0001001100001_1001110100110110100000_010011110110101110001010110011;
76 : data <= 65'b0001001011110_1001110110000010001110_010011110011101001101010000010;
77 : data <= 65'b0001001011010_1001110111001101011111_010011110000100101101110110111;
78 : data <= 65'b0001001010111_1001111000011000010011_010011101101100010011001000101;
79 : data <= 65'b0001001010011_1001111001100010101011_010011101010011111101000011100;
80 : data <= 65'b0001001010000_1001111010101100100111_010011100111011101011100101111;
81 : data <= 65'b0001001001100_1001111011110110000110_010011100100011011110101110000;
82 : data <= 65'b0001001001001_1001111100111111001011_010011100001011010110011010000;
83 : data <= 65'b0001001000101_1001111110000111110011_010011011110011010010101000011;
84 : data <= 65'b0001001000010_1001111111010000000001_010011011011011010011010111011;
85 : data <= 65'b0001000111110_1010000000010111110011_010011011000011011000100101001;
86 : data <= 65'b0001000111011_1010000001011111001011_010011010101011100010010000001;
87 : data <= 65'b0001000111000_1010000010100110001001_010011010010011110000010110110;
88 : data <= 65'b0001000110100_1010000011101100101100_010011001111100000010110111010;
89 : data <= 65'b0001000110001_1010000100110010110101_010011001100100011001110000001;
90 : data <= 65'b0001000101110_1010000101111000100100_010011001001100110100111111100;
91 : data <= 65'b0001000101011_1010000110111101111010_010011000110101010100100100001;
92 : data <= 65'b0001000101000_1010001000000010110111_010011000011101111000011100001;
93 : data <= 65'b0001000100100_1010001001000111011010_010011000000110100000100110001;
94 : data <= 65'b0001000100001_1010001010001011100100_010010111101111001101000000100;
95 : data <= 65'b0001000011110_1010001011001111010110_010010111010111111101101001101;
96 : data <= 65'b0001000011011_1010001100010010101111_010010111000000110010100000001;
97 : data <= 65'b0001000011000_1010001101010101110000_010010110101001101011100010011;
98 : data <= 65'b0001000010101_1010001110011000011000_010010110010010101000101110111;
99 : data <= 65'b0001000010010_1010001111011010101001_010010101111011101010000100001;
100 : data <= 65'b0001000001111_1010010000011100100010_010010101100100101111100000101;
101 : data <= 65'b0001000001100_1010010001011110000100_010010101001101111001000011000;
102 : data <= 65'b0001000001001_1010010010011111001110_010010100110111000110101001101;
103 : data <= 65'b0001000000110_1010010011100000000001_010010100100000011000010011010;
104 : data <= 65'b0001000000100_1010010100100000011110_010010100001001101101111110011;
105 : data <= 65'b0001000000001_1010010101100000100011_010010011110011000111101001100;
106 : data <= 65'b0000111111110_1010010110100000010010_010010011011100100101010011011;
107 : data <= 65'b0000111111011_1010010111011111101011_010010011000110000110111010100;
108 : data <= 65'b0000111111000_1010011000011110101110_010010010101111101100011101011;
109 : data <= 65'b0000111110110_1010011001011101011010_010010010011001010101111010111;
110 : data <= 65'b0000111110011_1010011010011011110001_010010010000011000011010001011;
111 : data <= 65'b0000111110000_1010011011011001110010_010010001101100110100011111110;
112 : data <= 65'b0000111101110_1010011100010111011110_010010001010110101001100100101;
113 : data <= 65'b0000111101011_1010011101010100110100_010010001000000100010011110100;
114 : data <= 65'b0000111101000_1010011110010001110101_010010000101010011111001100001;
115 : data <= 65'b0000111100110_1010011111001110100010_010010000010100011111101100011;
116 : data <= 65'b0000111100011_1010100000001010111001_010001111111110100011111101110;
117 : data <= 65'b0000111100000_1010100001000110111100_010001111101000101011111111000;
118 : data <= 65'b0000111011110_1010100010000010101011_010001111010010110111101110111;
119 : data <= 65'b0000111011011_1010100010111110000101_010001110111101000111001100000;
120 : data <= 65'b0000111011001_1010100011111001001011_010001110100111011010010101011;
121 : data <= 65'b0000111010110_1010100100110011111101_010001110010001110001001001100;
122 : data <= 65'b0000111010100_1010100101101110011011_010001101111100001011100111010;
123 : data <= 65'b0000111010001_1010100110101000100110_010001101100110101001101101011;
124 : data <= 65'b0000111001111_1010100111100010011101_010001101010001001011011010110;
125 : data <= 65'b0000111001101_1010101000011100000001_010001100111011110000101110000;
126 : data <= 65'b0000111001010_1010101001010101010010_010001100100110011001100110000;
127 : data <= 65'b0000111001000_1010101010001110010000_010001100010001000110000001100;
128 : data <= 65'b0000111000101_1010101011000110111010_010001011111011110101111111100;
129 : data <= 65'b0000111000011_1010101011111111010010_010001011100110101001011110101;
130 : data <= 65'b0000111000001_1010101100110111011000_010001011010001100000011101110;
131 : data <= 65'b0000110111110_1010101101101111001011_010001010111100011010111011111;
132 : data <= 65'b0000110111100_1010101110100110101011_010001010100111011000110111110;
133 : data <= 65'b0000110111010_1010101111011101111010_010001010010010011010010000001;
134 : data <= 65'b0000110111000_1010110000010100110110_010001001111101011111000100001;
135 : data <= 65'b0000110110101_1010110001001011100001_010001001101000100111010010011;
136 : data <= 65'b0000110110011_1010110010000001111010_010001001010011110010111010000;
137 : data <= 65'b0000110110001_1010110010111000000001_010001000111111000001111001110;
138 : data <= 65'b0000110101111_1010110011101101110110_010001000101010010100010000100;
139 : data <= 65'b0000110101101_1010110100100011011011_010001000010101101001111101010;
140 : data <= 65'b0000110101010_1010110101011000101110_010001000000001000010111110111;
141 : data <= 65'b0000110101000_1010110110001101110000_010000111101100011111010100011;
142 : data <= 65'b0000110100110_1010110111000010100001_010000111010111111110111100110;
143 : data <= 65'b0000110100100_1010110111110111000001_010000111000011100001110110110;
144 : data <= 65'b0000110100010_1010111000101011010000_010000110101111001000000001011;
145 : data <= 65'b0000110100000_1010111001011111001111_010000110011010110001011011101;
146 : data <= 65'b0000110011110_1010111010010010111110_010000110000110011110000100101;
147 : data <= 65'b0000110011100_1010111011000110011100_010000101110010001101111011001;
148 : data <= 65'b0000110011010_1010111011111001101010_010000101011110000000111110001;
149 : data <= 65'b0000110011000_1010111100101100100111_010000101001001110111001100111;
150 : data <= 65'b0000110010110_1010111101011111010101_010000100110101110000100110000;
151 : data <= 65'b0000110010100_1010111110010001110011_010000100100001101101001000111;
152 : data <= 65'b0000110010010_1010111111000100000001_010000100001101101100110100010;
153 : data <= 65'b0000110010000_1010111111110101111111_010000011111001101111100111010;
154 : data <= 65'b0000110001110_1011000000100111101110_010000011100101110101100000111;
155 : data <= 65'b0000110001100_1011000001011001001110_010000011010001111110100000001;
156 : data <= 65'b0000110001010_1011000010001010011110_010000010111110001010100100010;
157 : data <= 65'b0000110001000_1011000010111011011111_010000010101010011001101100000;
158 : data <= 65'b0000110000110_1011000011101100010001_010000010010110101011110110110;
159 : data <= 65'b0000110000100_1011000100011100110100_010000010000011000001000011010;
160 : data <= 65'b0000110000011_1011000101001101001000_010000001101111011001010000110;
161 : data <= 65'b0000110000001_1011000101111101001101_010000001011011110100011110011;
162 : data <= 65'b0000101111111_1011000110101101000100_010000001001000010010101011001;
163 : data <= 65'b0000101111101_1011000111011100101100_010000000110100110011110110000;
164 : data <= 65'b0000101111011_1011001000001100000110_010000000100001010111111110010;
165 : data <= 65'b0000101111001_1011001000111011010001_010000000001101111111000010111;
166 : data <= 65'b0000101111000_1011001001101010001110_001111111111010101001000011001;
167 : data <= 65'b0000101110110_1011001010011000111101_001111111100111010101111110000;
168 : data <= 65'b0000101110100_1011001011000111011110_001111111010100000101110010101;
169 : data <= 65'b0000101110010_1011001011110101110001_001111111000000111000100000001;
170 : data <= 65'b0000101110001_1011001100100011110110_001111110101101101110000101110;
171 : data <= 65'b0000101101111_1011001101010001101110_001111110011010100110100010100;
172 : data <= 65'b0000101101101_1011001101111111011000_001111110000111100001110101100;
173 : data <= 65'b0000101101100_1011001110101100110100_001111101110100011111111110000;
174 : data <= 65'b0000101101010_1011001111011010000010_001111101100001100000111011010;
175 : data <= 65'b0000101101000_1011010000000111000100_001111101001110100100101100010;
176 : data <= 65'b0000101100111_1011010000110011111000_001111100111011101011010000001;
177 : data <= 65'b0000101100101_1011010001100000011111_001111100101000110100100110010;
178 : data <= 65'b0000101100011_1011010010001100111001_001111100010110000000101101101;
179 : data <= 65'b0000101100010_1011010010111001000101_001111100000011001111100101101;
180 : data <= 65'b0000101100000_1011010011100101000101_001111011110000100001001101010;
181 : data <= 65'b0000101011110_1011010100010000111000_001111011011101110101100011111;
182 : data <= 65'b0000101011101_1011010100111100011110_001111011001011001100101000100;
183 : data <= 65'b0000101011011_1011010101100111111000_001111010111000100110011010100;
184 : data <= 65'b0000101011010_1011010110010011000101_001111010100110000010111001000;
185 : data <= 65'b0000101011000_1011010110111110000110_001111010010011100010000011011;
186 : data <= 65'b0000101010111_1011010111101000111010_001111010000001000011111000101;
187 : data <= 65'b0000101010101_1011011000010011100010_001111001101110101000011000001;
188 : data <= 65'b0000101010100_1011011000111101111101_001111001011100001111100001000;
189 : data <= 65'b0000101010010_1011011001101000001101_001111001001001111001010010101;
190 : data <= 65'b0000101010000_1011011010010010010000_001111000110111100101101100010;
191 : data <= 65'b0000101001111_1011011010111100001000_001111000100101010100101101000;
192 : data <= 65'b0000101001101_1011011011100101110011_001111000010011000110010100001;
193 : data <= 65'b0000101001100_1011011100001111010011_001111000000000111010100001000;
194 : data <= 65'b0000101001011_1011011100111000100111_001110111101110110001010010111;
195 : data <= 65'b0000101001001_1011011101100001101111_001110111011100101010101001000;
196 : data <= 65'b0000101001000_1011011110001010101100_001110111001010100110100010101;
197 : data <= 65'b0000101000110_1011011110110011011101_001110110111000100100111111001;
198 : data <= 65'b0000101000101_1011011111011100000011_001110110100110100101111101101;
199 : data <= 65'b0000101000011_1011100000000100011101_001110110010100101001011101100;
200 : data <= 65'b0000101000010_1011100000101100101100_001110110000010101111011110000;
201 : data <= 65'b0000101000001_1011100001010100110000_001110101110000110111111110100;
202 : data <= 65'b0000100111111_1011100001111100101000_001110101011111000010111110010;
203 : data <= 65'b0000100111110_1011100010100100010110_001110101001101010000011100101;
204 : data <= 65'b0000100111100_1011100011001011111001_001110100111011100000011000111;
205 : data <= 65'b0000100111011_1011100011110011010000_001110100101001110010110010011;
206 : data <= 65'b0000100111010_1011100100011010011101_001110100011000000111101000010;
207 : data <= 65'b0000100111000_1011100101000001011111_001110100000110011110111010001;
208 : data <= 65'b0000100110111_1011100101101000010110_001110011110100111000100111001;
209 : data <= 65'b0000100110110_1011100110001111000011_001110011100011010100101110110;
210 : data <= 65'b0000100110100_1011100110110101100101_001110011010001110011010000001;
211 : data <= 65'b0000100110011_1011100111011011111101_001110011000000010100001010110;
212 : data <= 65'b0000100110010_1011101000000010001010_001110010101110110111011101111;
213 : data <= 65'b0000100110000_1011101000101000001100_001110010011101011101001001000;
214 : data <= 65'b0000100101111_1011101001001110000101_001110010001100000101001011010;
215 : data <= 65'b0000100101110_1011101001110011110011_001110001111010101111100100001;
216 : data <= 65'b0000100101101_1011101010011001010111_001110001101001011100010011001;
217 : data <= 65'b0000100101011_1011101010111110110001_001110001011000001011010111011;
218 : data <= 65'b0000100101010_1011101011100100000001_001110001000110111100110000011;
219 : data <= 65'b0000100101001_1011101100001001000110_001110000110101110000011101011;
220 : data <= 65'b0000100101000_1011101100101110000010_001110000100100100110011110000;
221 : data <= 65'b0000100100110_1011101101010010110100_001110000010011011110110001011;
222 : data <= 65'b0000100100101_1011101101110111011100_001110000000010011001010111000;
223 : data <= 65'b0000100100100_1011101110011011111011_001101111110001010110001110011;
224 : data <= 65'b0000100100011_1011101111000000001111_001101111100000010101010110101;
225 : data <= 65'b0000100100001_1011101111100100011011_001101111001111010110101111011;
226 : data <= 65'b0000100100000_1011110000001000011100_001101110111110011010011000000;
227 : data <= 65'b0000100011111_1011110000101100010100_001101110101101100000001111111;
228 : data <= 65'b0000100011110_1011110001010000000011_001101110011100101000010110011;
229 : data <= 65'b0000100011101_1011110001110011101000_001101110001011110010101010111;
230 : data <= 65'b0000100011100_1011110010010111000100_001101101111010111111001101000;
231 : data <= 65'b0000100011010_1011110010111010010110_001101101101010001101111011111;
232 : data <= 65'b0000100011001_1011110011011101100000_001101101011001011110110111001;
233 : data <= 65'b0000100011000_1011110100000000100000_001101101001000110001111110001;
234 : data <= 65'b0000100010111_1011110100100011010111_001101100111000000111010000011;
235 : data <= 65'b0000100010110_1011110101000110000101_001101100100111011110101101001;
236 : data <= 65'b0000100010101_1011110101101000101010_001101100010110111000010100000;
237 : data <= 65'b0000100010100_1011110110001011000110_001101100000110010100000100100;
238 : data <= 65'b0000100010010_1011110110101101011001_001101011110101110001111101110;
239 : data <= 65'b0000100010001_1011110111001111100100_001101011100101010001111111100;
240 : data <= 65'b0000100010000_1011110111110001100101_001101011010100110100001001000;
241 : data <= 65'b0000100001111_1011111000010011011110_001101011000100011000011001111;
242 : data <= 65'b0000100001110_1011111000110101001111_001101010110011111110110001100;
243 : data <= 65'b0000100001101_1011111001010110110110_001101010100011100111001111011;
244 : data <= 65'b0000100001100_1011111001111000010101_001101010010011010001110010111;
245 : data <= 65'b0000100001011_1011111010011001101100_001101010000010111110011011101;
246 : data <= 65'b0000100001010_1011111010111010111010_001101001110010101101001000111;
247 : data <= 65'b0000100001001_1011111011011011111111_001101001100010011101111010010;
248 : data <= 65'b0000100001000_1011111011111100111100_001101001010010010000101111010;
249 : data <= 65'b0000100000111_1011111100011101110001_001101001000010000101100111010;
250 : data <= 65'b0000100000110_1011111100111110011110_001101000110001111100100001111;
251 : data <= 65'b0000100000101_1011111101011111000010_001101000100001110101011110100;
252 : data <= 65'b0000100000100_1011111101111111011111_001101000010001110000011100101;
253 : data <= 65'b0000100000011_1011111110011111110011_001101000000001101101011011110;
254 : data <= 65'b0000100000010_1011111110111111111111_001100111110001101100011011011;
255 : data <= 65'b0000100000000_1011111111100000000011_001100111100001101101011011000;
endcase
end

endmodule
