//Table with Sqrt2 Coefficient values

module Sqrt2_Coeffs (
clk,     // Clock
address, // Address input
data    // Data output
);
input clk;
input [5:0] address;
output [31:0] data;
reg [31:0] data ;
       
always@(clk)
begin
case(address)
0 : data = 32'b00000000001111111100_010000000000;	
1 : data = 32'b00000000001111110100_010111111010;
2 : data = 32'b00000000001111101100_011111101100;
3 : data = 32'b00000000001111100101_000111011000;			//Coefficient values
4 : data = 32'b00000000001111011101_001110111100;
5 : data = 32'b00000000001111010110_010110011001;
6 : data = 32'b00000000001111001111_011101110000;
7 : data = 32'b00000000001111001000_000101000000;
8 : data = 32'b00000000001111000010_001100001010;
9 : data = 32'b00000000001110111011_010011001110;
10 : data = 32'b00000000001110110101_011010001100;
11 : data = 32'b00000000001110101110_000001000100;
12 : data = 32'b00000000001110101000_000111110111;
13 : data = 32'b00000000001110100010_001110100101;
14 : data = 32'b00000000001110011100_010101001101;
15 : data = 32'b00000000001110010110_011011110000;
16 : data = 32'b00000000001110010001_000010001111;
17 : data = 32'b00000000001110001011_001000101000;
18 : data = 32'b00000000001110000101_001110111101;
19 : data = 32'b00000000001110000000_010101001101;
20 : data = 32'b00000000001101111011_011011011001;
21 : data = 32'b00000000001101110101_000001100001;
22 : data = 32'b00000000001101110000_000111100100;
23 : data = 32'b00000000001101101011_001101100011;
24 : data = 32'b00000000001101100110_010011011111;
25 : data = 32'b00000000001101100001_011001010110;
26 : data = 32'b00000000001101011101_011111001010;
27 : data = 32'b00000000001101011000_000100111001;
28 : data = 32'b00000000001101010011_001010100110;
29 : data = 32'b00000000001101001111_010000001110;
30 : data = 32'b00000000001101001010_010101110100;
31 : data = 32'b00000000001101000110_011011010101;
32 : data = 32'b00000000001101000001_000000110100;
33 : data = 32'b00000000001100111101_000110001111;
34 : data = 32'b00000000001100111001_001011100111;
35 : data = 32'b00000000001100110101_010000111101;
36 : data = 32'b00000000001100110001_010110001111;
37 : data = 32'b00000000001100101101_011011011110;
38 : data = 32'b00000000001100101001_000000101010;
39 : data = 32'b00000000001100100101_000101110011;
40 : data = 32'b00000000001100100001_001010111010;
41 : data = 32'b00000000001100011101_001111111110;
42 : data = 32'b00000000001100011001_010100111111;
43 : data = 32'b00000000001100010110_011001111101;
44 : data = 32'b00000000001100010010_011110111001;
45 : data = 32'b00000000001100001110_000011110011;
46 : data = 32'b00000000001100001011_001000101010;
47 : data = 32'b00000000001100000111_001101011111;
48 : data = 32'b00000000001100000100_010010010001;
49 : data = 32'b00000000001100000000_010111000001;
50 : data = 32'b00000000001011111101_011011101111;
51 : data = 32'b00000000001011111010_000000011010;
52 : data = 32'b00000000001011110110_000101000011;
53 : data = 32'b00000000001011110011_001001101010;
54 : data = 32'b00000000001011110000_001110001111;
55 : data = 32'b00000000001011101101_010010110010;
56 : data = 32'b00000000001011101010_010111010011;
57 : data = 32'b00000000001011100111_011011110010;
58 : data = 32'b00000000001011100100_000000001110;
59 : data = 32'b00000000001011100001_000100101001;
60 : data = 32'b00000000001011011110_001001000010;
61 : data = 32'b00000000001011011011_001101011001;
62 : data = 32'b00000000001011011000_010001101111;
63 : data = 32'b00000000001011010101_010110000010;
endcase
end

endmodule
